module window_processor_top (
    data_in,
    row_size,
    data_in_valid,
    enable,
    clear,
    clock,
    col_size,
    start,
    data_out,
    data_out_valid,
    idle,
    last_in,
    last_out,
    ready,
    total_count
);

    input [15:0] data_in;
    input [9:0] row_size;
    input data_in_valid;
    input enable;
    input clear;
    input clock;
    input [9:0] col_size;
    input start;
    output [15:0] data_out;
    output data_out_valid;
    output idle;
    output last_in;
    output last_out;
    output ready;
    output [20:0] total_count;

    wire [20:0] _84;
    wire [20:0] _160;
    wire [20:0] _156;
    wire [20:0] _157;
    wire _146;
    wire [3:0] _145;
    wire [4:0] _147;
    wire _143;
    wire [4:0] _144;
    wire [4:0] _148;
    wire _139;
    wire [4:0] _140;
    wire _136;
    wire [4:0] _137;
    wire [4:0] _141;
    wire [4:0] _149;
    wire _131;
    wire [4:0] _132;
    wire _128;
    wire [4:0] _129;
    wire [4:0] _133;
    wire _124;
    wire [4:0] _125;
    wire _121;
    wire [4:0] _122;
    wire [4:0] _126;
    wire [4:0] _134;
    wire [4:0] _150;
    wire _115;
    wire [4:0] _116;
    wire _112;
    wire [4:0] _113;
    wire [4:0] _117;
    wire _108;
    wire [4:0] _109;
    wire _105;
    wire [4:0] _106;
    wire [4:0] _110;
    wire [4:0] _118;
    wire _100;
    wire [4:0] _101;
    wire _97;
    wire [4:0] _98;
    wire [4:0] _102;
    wire _93;
    wire [4:0] _94;
    wire [15:0] _1;
    wire [15:0] _88;
    wire [15:0] _72;
    reg [15:0] _73;
    wire [15:0] o$result$prev;
    wire [15:0] _3;
    wire [15:0] _89;
    wire _90;
    wire [4:0] _91;
    wire [4:0] _95;
    wire [4:0] _103;
    wire [4:0] _119;
    wire [4:0] _151;
    wire [20:0] _152;
    wire [20:0] _153;
    wire _4;
    wire [20:0] _154;
    wire _82;
    wire [20:0] _155;
    wire _80;
    wire [20:0] _158;
    wire _78;
    wire [20:0] _161;
    wire [20:0] _5;
    reg [20:0] _85;
    wire [20:0] o$total_count;
    wire _162;
    wire _165;
    wire o$ready;
    wire _171;
    reg _170;
    wire _172;
    wire o$last_out;
    wire o$last_in;
    wire o$idle;
    wire i$data_in$valid1;
    reg _226;
    reg _229;
    reg _232;
    wire o$result$valid;
    reg _235;
    wire _237;
    wire o$data_out_valid;
    wire [3:0] _1013;
    wire _1008;
    wire [2:0] _1007;
    wire [3:0] _1009;
    wire _1005;
    wire [3:0] _1006;
    wire [3:0] _1010;
    wire _1001;
    wire [3:0] _1002;
    wire _998;
    wire [3:0] _999;
    wire [3:0] _1003;
    wire [3:0] _1011;
    wire _993;
    wire [3:0] _994;
    wire _990;
    wire [3:0] _991;
    wire [3:0] _995;
    wire _986;
    wire [3:0] _987;
    wire _981;
    wire _980;
    wire _979;
    wire _978;
    wire _977;
    wire _976;
    wire _975;
    wire _974;
    wire [7:0] _982;
    wire _983;
    wire [3:0] _984;
    wire [3:0] _988;
    wire [3:0] _996;
    wire [3:0] _1012;
    wire _1014;
    wire _966;
    wire [3:0] _967;
    wire _963;
    wire [3:0] _964;
    wire [3:0] _968;
    wire _959;
    wire [3:0] _960;
    wire _956;
    wire [3:0] _957;
    wire [3:0] _961;
    wire [3:0] _969;
    wire _951;
    wire [3:0] _952;
    wire _948;
    wire [3:0] _949;
    wire [3:0] _953;
    wire _944;
    wire [3:0] _945;
    wire _939;
    wire _938;
    wire _937;
    wire _936;
    wire _935;
    wire _934;
    wire _933;
    wire _932;
    wire [7:0] _940;
    wire _941;
    wire [3:0] _942;
    wire [3:0] _946;
    wire [3:0] _954;
    wire [3:0] _970;
    wire _972;
    wire _924;
    wire [3:0] _925;
    wire _921;
    wire [3:0] _922;
    wire [3:0] _926;
    wire _917;
    wire [3:0] _918;
    wire _914;
    wire [3:0] _915;
    wire [3:0] _919;
    wire [3:0] _927;
    wire _909;
    wire [3:0] _910;
    wire _906;
    wire [3:0] _907;
    wire [3:0] _911;
    wire _902;
    wire [3:0] _903;
    wire _897;
    wire _896;
    wire _895;
    wire _894;
    wire _893;
    wire _892;
    wire _891;
    wire _890;
    wire [7:0] _898;
    wire _899;
    wire [3:0] _900;
    wire [3:0] _904;
    wire [3:0] _912;
    wire [3:0] _928;
    wire _930;
    wire _882;
    wire [3:0] _883;
    wire _879;
    wire [3:0] _880;
    wire [3:0] _884;
    wire _875;
    wire [3:0] _876;
    wire _872;
    wire [3:0] _873;
    wire [3:0] _877;
    wire [3:0] _885;
    wire _867;
    wire [3:0] _868;
    wire _864;
    wire [3:0] _865;
    wire [3:0] _869;
    wire _860;
    wire [3:0] _861;
    wire _855;
    wire _854;
    wire _853;
    wire _852;
    wire _851;
    wire _850;
    wire _849;
    wire _848;
    wire [7:0] _856;
    wire _857;
    wire [3:0] _858;
    wire [3:0] _862;
    wire [3:0] _870;
    wire [3:0] _886;
    wire _888;
    wire _840;
    wire [3:0] _841;
    wire _837;
    wire [3:0] _838;
    wire [3:0] _842;
    wire _833;
    wire [3:0] _834;
    wire _830;
    wire [3:0] _831;
    wire [3:0] _835;
    wire [3:0] _843;
    wire _825;
    wire [3:0] _826;
    wire _822;
    wire [3:0] _823;
    wire [3:0] _827;
    wire _818;
    wire [3:0] _819;
    wire _813;
    wire _812;
    wire _811;
    wire _810;
    wire _809;
    wire _808;
    wire _807;
    wire _806;
    wire [7:0] _814;
    wire _815;
    wire [3:0] _816;
    wire [3:0] _820;
    wire [3:0] _828;
    wire [3:0] _844;
    wire _846;
    wire _798;
    wire [3:0] _799;
    wire _795;
    wire [3:0] _796;
    wire [3:0] _800;
    wire _791;
    wire [3:0] _792;
    wire _788;
    wire [3:0] _789;
    wire [3:0] _793;
    wire [3:0] _801;
    wire _783;
    wire [3:0] _784;
    wire _780;
    wire [3:0] _781;
    wire [3:0] _785;
    wire _776;
    wire [3:0] _777;
    wire _771;
    wire _770;
    wire _769;
    wire _768;
    wire _767;
    wire _766;
    wire _765;
    wire _764;
    wire [7:0] _772;
    wire _773;
    wire [3:0] _774;
    wire [3:0] _778;
    wire [3:0] _786;
    wire [3:0] _802;
    wire _804;
    wire _756;
    wire [3:0] _757;
    wire _753;
    wire [3:0] _754;
    wire [3:0] _758;
    wire _749;
    wire [3:0] _750;
    wire _746;
    wire [3:0] _747;
    wire [3:0] _751;
    wire [3:0] _759;
    wire _741;
    wire [3:0] _742;
    wire _738;
    wire [3:0] _739;
    wire [3:0] _743;
    wire _734;
    wire [3:0] _735;
    wire _729;
    wire _728;
    wire _727;
    wire _726;
    wire _725;
    wire _724;
    wire _723;
    wire _722;
    wire [7:0] _730;
    wire _731;
    wire [3:0] _732;
    wire [3:0] _736;
    wire [3:0] _744;
    wire [3:0] _760;
    wire _762;
    wire _714;
    wire [3:0] _715;
    wire _711;
    wire [3:0] _712;
    wire [3:0] _716;
    wire _707;
    wire [3:0] _708;
    wire _704;
    wire [3:0] _705;
    wire [3:0] _709;
    wire [3:0] _717;
    wire _699;
    wire [3:0] _700;
    wire _696;
    wire [3:0] _697;
    wire [3:0] _701;
    wire _692;
    wire [3:0] _693;
    wire _687;
    wire _686;
    wire _685;
    wire _684;
    wire _683;
    wire _682;
    wire _681;
    wire _680;
    wire [7:0] _688;
    wire _689;
    wire [3:0] _690;
    wire [3:0] _694;
    wire [3:0] _702;
    wire [3:0] _718;
    wire _720;
    wire _672;
    wire [3:0] _673;
    wire _669;
    wire [3:0] _670;
    wire [3:0] _674;
    wire _665;
    wire [3:0] _666;
    wire _662;
    wire [3:0] _663;
    wire [3:0] _667;
    wire [3:0] _675;
    wire _657;
    wire [3:0] _658;
    wire _654;
    wire [3:0] _655;
    wire [3:0] _659;
    wire _650;
    wire [3:0] _651;
    wire _645;
    wire _644;
    wire _643;
    wire _642;
    wire _641;
    wire _640;
    wire _639;
    wire _638;
    wire [7:0] _646;
    wire _647;
    wire [3:0] _648;
    wire [3:0] _652;
    wire [3:0] _660;
    wire [3:0] _676;
    wire _678;
    wire _630;
    wire [3:0] _631;
    wire _627;
    wire [3:0] _628;
    wire [3:0] _632;
    wire _623;
    wire [3:0] _624;
    wire _620;
    wire [3:0] _621;
    wire [3:0] _625;
    wire [3:0] _633;
    wire _615;
    wire [3:0] _616;
    wire _612;
    wire [3:0] _613;
    wire [3:0] _617;
    wire _608;
    wire [3:0] _609;
    wire _603;
    wire _602;
    wire _601;
    wire _600;
    wire _599;
    wire _598;
    wire _597;
    wire _596;
    wire [7:0] _604;
    wire _605;
    wire [3:0] _606;
    wire [3:0] _610;
    wire [3:0] _618;
    wire [3:0] _634;
    wire _636;
    wire _588;
    wire [3:0] _589;
    wire _585;
    wire [3:0] _586;
    wire [3:0] _590;
    wire _581;
    wire [3:0] _582;
    wire _578;
    wire [3:0] _579;
    wire [3:0] _583;
    wire [3:0] _591;
    wire _573;
    wire [3:0] _574;
    wire _570;
    wire [3:0] _571;
    wire [3:0] _575;
    wire _566;
    wire [3:0] _567;
    wire _561;
    wire _560;
    wire _559;
    wire _558;
    wire _557;
    wire _556;
    wire _555;
    wire _554;
    wire [7:0] _562;
    wire _563;
    wire [3:0] _564;
    wire [3:0] _568;
    wire [3:0] _576;
    wire [3:0] _592;
    wire _594;
    wire _546;
    wire [3:0] _547;
    wire _543;
    wire [3:0] _544;
    wire [3:0] _548;
    wire _539;
    wire [3:0] _540;
    wire _536;
    wire [3:0] _537;
    wire [3:0] _541;
    wire [3:0] _549;
    wire _531;
    wire [3:0] _532;
    wire _528;
    wire [3:0] _529;
    wire [3:0] _533;
    wire _524;
    wire [3:0] _525;
    wire _519;
    wire _518;
    wire _517;
    wire _516;
    wire _515;
    wire _514;
    wire _513;
    wire _512;
    wire [7:0] _520;
    wire _521;
    wire [3:0] _522;
    wire [3:0] _526;
    wire [3:0] _534;
    wire [3:0] _550;
    wire _552;
    wire _504;
    wire [3:0] _505;
    wire _501;
    wire [3:0] _502;
    wire [3:0] _506;
    wire _497;
    wire [3:0] _498;
    wire _494;
    wire [3:0] _495;
    wire [3:0] _499;
    wire [3:0] _507;
    wire _489;
    wire [3:0] _490;
    wire _486;
    wire [3:0] _487;
    wire [3:0] _491;
    wire _482;
    wire [3:0] _483;
    wire _477;
    wire _476;
    wire _475;
    wire _474;
    wire _473;
    wire _472;
    wire _471;
    wire _470;
    wire [7:0] _478;
    wire _479;
    wire [3:0] _480;
    wire [3:0] _484;
    wire [3:0] _492;
    wire [3:0] _508;
    wire _510;
    wire _462;
    wire [3:0] _463;
    wire _459;
    wire [3:0] _460;
    wire [3:0] _464;
    wire _455;
    wire [3:0] _456;
    wire _452;
    wire [3:0] _453;
    wire [3:0] _457;
    wire [3:0] _465;
    wire _447;
    wire [3:0] _448;
    wire _444;
    wire [3:0] _445;
    wire [3:0] _449;
    wire _440;
    wire [3:0] _441;
    wire _435;
    wire _434;
    wire _433;
    wire _432;
    wire _431;
    wire _430;
    wire _429;
    wire _428;
    wire [7:0] _436;
    wire _437;
    wire [3:0] _438;
    wire [3:0] _442;
    wire [3:0] _450;
    wire [3:0] _466;
    wire _468;
    wire _420;
    wire [3:0] _421;
    wire _417;
    wire [3:0] _418;
    wire [3:0] _422;
    wire _413;
    wire [3:0] _414;
    wire _410;
    wire [3:0] _411;
    wire [3:0] _415;
    wire [3:0] _423;
    wire _405;
    wire [3:0] _406;
    wire _402;
    wire [3:0] _403;
    wire [3:0] _407;
    wire _398;
    wire [3:0] _399;
    wire _393;
    wire _392;
    wire _391;
    wire _390;
    wire _389;
    wire _388;
    wire _387;
    wire _386;
    wire [7:0] _394;
    wire _395;
    wire [3:0] _396;
    wire [3:0] _400;
    wire [3:0] _408;
    wire [3:0] _424;
    wire _426;
    wire _378;
    wire [3:0] _379;
    wire _375;
    wire [3:0] _376;
    wire [3:0] _380;
    wire _371;
    wire [3:0] _372;
    wire _368;
    wire [3:0] _369;
    wire [3:0] _373;
    wire [3:0] _381;
    wire _363;
    wire [3:0] _364;
    wire _360;
    wire [3:0] _361;
    wire [3:0] _365;
    wire _356;
    wire [3:0] _357;
    wire [46:0] _347;
    wire [47:0] _349;
    wire [15:0] _350;
    wire _351;
    wire [15:0] _345;
    wire _346;
    wire [15:0] _338;
    wire [15:0] _339;
    wire [15:0] _337;
    wire [15:0] i$data_in$d2;
    reg [15:0] _329;
    reg [15:0] _332;
    reg [15:0] _335;
    wire i$data_in$bottom1;
    reg _321;
    reg _324;
    wire [15:0] _325;
    wire [15:0] _326;
    wire [15:0] _336;
    wire [47:0] _340;
    wire [46:0] _341;
    wire [47:0] _342;
    wire [15:0] _343;
    wire _344;
    wire [46:0] _313;
    wire [47:0] _315;
    wire [15:0] _316;
    wire _317;
    wire [15:0] _307;
    reg [15:0] _305;
    wire [15:0] _306;
    wire [47:0] _308;
    wire [46:0] _309;
    wire [47:0] _310;
    wire [15:0] _311;
    wire _312;
    wire [46:0] _297;
    wire [47:0] _299;
    wire [15:0] _300;
    wire _301;
    wire [15:0] _295;
    wire _296;
    wire i$data_in$right1;
    reg _283;
    reg _286;
    wire [15:0] _287;
    wire [15:0] _288;
    wire [15:0] _289;
    wire [15:0] _280;
    wire _223;
    wire _238;
    wire _239;
    wire [21:0] _247;
    reg [21:0] _248[0:1023];
    wire [9:0] _241;
    reg [9:0] _242;
    wire [21:0] _249;
    wire [15:0] _250;
    wire [15:0] i$data_in$d0;
    reg [15:0] _272;
    reg [15:0] _275;
    reg [15:0] _278;
    wire _243;
    wire i$data_in$left1;
    reg _264;
    reg _267;
    wire [15:0] _268;
    wire [15:0] _259;
    wire _244;
    wire i$data_in$top1;
    reg _255;
    reg _258;
    wire [15:0] _261;
    wire [15:0] _269;
    wire [15:0] _279;
    wire [47:0] _290;
    wire [46:0] _291;
    wire [47:0] _292;
    wire [15:0] _293;
    wire _294;
    wire [7:0] _352;
    wire _353;
    wire [3:0] _354;
    wire [3:0] _358;
    wire [3:0] _366;
    wire [3:0] _382;
    wire _384;
    wire [15:0] _1015;
    wire [15:0] _1016;
    wire [15:0] _246;
    wire [15:0] i$data_in$d1;
    reg [15:0] _67;
    reg [15:0] _70;
    wire [15:0] _1017;
    reg [15:0] _1020;
    wire [15:0] o$result$d;
    reg [15:0] _1079;
    wire vdd;
    wire gnd;
    wire [1:0] _75;
    wire [1:0] _1075;
    wire [1:0] _1072;
    wire [1:0] _1073;
    wire i$enable;
    wire i$clear;
    wire i$clock;
    wire _218;
    wire _217;
    wire _219;
    wire _220;
    wire [15:0] _32;
    wire [15:0] i$data_in;
    wire [9:0] _185;
    wire [9:0] _186;
    wire _190;
    wire [9:0] _177;
    wire _181;
    wire _191;
    wire _215;
    wire [9:0] _35;
    wire [9:0] i$row_size;
    wire [9:0] _1022;
    wire _1021;
    wire [9:0] _1023;
    wire [9:0] _37;
    reg [9:0] _180;
    wire [9:0] _1038;
    wire [9:0] _1034;
    wire [9:0] _1035;
    wire [9:0] _1031;
    wire [9:0] _1032;
    wire _1026;
    wire [9:0] _1033;
    wire _1025;
    wire [9:0] _1036;
    wire _1024;
    wire [9:0] _1039;
    wire [9:0] _38;
    reg [9:0] _175;
    wire [9:0] _212;
    wire _213;
    wire _210;
    wire [9:0] _207;
    wire _208;
    wire [21:0] _216;
    reg [21:0] _221[0:1023];
    wire _202;
    wire _201;
    wire _203;
    wire _204;
    wire [9:0] _197;
    wire [9:0] _1053;
    wire [9:0] _1049;
    wire _40;
    wire i$data_in_valid;
    wire [9:0] _1050;
    wire _43;
    wire i$enable_0;
    wire _46;
    wire i$clear_0;
    wire _49;
    wire i$clock_0;
    wire [9:0] _52;
    wire [9:0] i$col_size;
    wire _55;
    wire i$start;
    wire [9:0] _1041;
    wire _1040;
    wire [9:0] _1042;
    wire [9:0] _57;
    reg [9:0] _189;
    wire [9:0] _1028;
    wire _1029;
    wire [9:0] _1047;
    wire _1045;
    wire [9:0] _1048;
    wire _1044;
    wire [9:0] _1051;
    wire _1043;
    wire [9:0] _1054;
    wire [9:0] _58;
    reg [9:0] _184;
    wire [9:0] _193;
    wire _194;
    wire [9:0] _198;
    reg [9:0] _205;
    wire [21:0] _222;
    wire _245;
    wire i$data_in$last1;
    reg _1057;
    reg _1060;
    reg _1063;
    wire o$result$last;
    wire _61;
    wire [1:0] _1070;
    wire [1:0] _1067;
    wire _1068;
    wire [1:0] _1069;
    wire [1:0] _81;
    wire _1066;
    wire [1:0] _1071;
    wire [1:0] _79;
    wire _1065;
    wire [1:0] _1074;
    wire _1064;
    wire [1:0] _1076;
    wire [1:0] _62;
    reg [1:0] _76;
    wire _166;
    wire _167;
    wire [15:0] _1081;
    wire [15:0] o$data_out;
    assign _84 = 21'b000000000000000000000;
    assign _160 = i$start ? _84 : _85;
    assign _156 = _4 ? _153 : _85;
    assign _157 = i$data_in_valid ? _156 : _85;
    assign _146 = _89[0:0];
    assign _145 = 4'b0000;
    assign _147 = { _145,
                    _146 };
    assign _143 = _89[1:1];
    assign _144 = { _145,
                    _143 };
    assign _148 = _144 + _147;
    assign _139 = _89[2:2];
    assign _140 = { _145,
                    _139 };
    assign _136 = _89[3:3];
    assign _137 = { _145,
                    _136 };
    assign _141 = _137 + _140;
    assign _149 = _141 + _148;
    assign _131 = _89[4:4];
    assign _132 = { _145,
                    _131 };
    assign _128 = _89[5:5];
    assign _129 = { _145,
                    _128 };
    assign _133 = _129 + _132;
    assign _124 = _89[6:6];
    assign _125 = { _145,
                    _124 };
    assign _121 = _89[7:7];
    assign _122 = { _145,
                    _121 };
    assign _126 = _122 + _125;
    assign _134 = _126 + _133;
    assign _150 = _134 + _149;
    assign _115 = _89[8:8];
    assign _116 = { _145,
                    _115 };
    assign _112 = _89[9:9];
    assign _113 = { _145,
                    _112 };
    assign _117 = _113 + _116;
    assign _108 = _89[10:10];
    assign _109 = { _145,
                    _108 };
    assign _105 = _89[11:11];
    assign _106 = { _145,
                    _105 };
    assign _110 = _106 + _109;
    assign _118 = _110 + _117;
    assign _100 = _89[12:12];
    assign _101 = { _145,
                    _100 };
    assign _97 = _89[13:13];
    assign _98 = { _145,
                   _97 };
    assign _102 = _98 + _101;
    assign _93 = _89[14:14];
    assign _94 = { _145,
                   _93 };
    assign _1 = o$result$d;
    assign _88 = ~ _1;
    assign _72 = 16'b0000000000000000;
    always @(posedge i$clock) begin
        if (i$clear)
            _73 <= _72;
        else
            if (i$enable)
                _73 <= _70;
    end
    assign o$result$prev = _73;
    assign _3 = o$result$prev;
    assign _89 = _3 & _88;
    assign _90 = _89[15:15];
    assign _91 = { _145,
                   _90 };
    assign _95 = _91 + _94;
    assign _103 = _95 + _102;
    assign _119 = _103 + _118;
    assign _151 = _119 + _150;
    assign _152 = { _72,
                    _151 };
    assign _153 = _85 + _152;
    assign _4 = o$result$valid;
    assign _154 = _4 ? _153 : _85;
    assign _82 = _76 == _81;
    assign _155 = _82 ? _154 : _85;
    assign _80 = _76 == _79;
    assign _158 = _80 ? _157 : _155;
    assign _78 = _76 == _75;
    assign _161 = _78 ? _160 : _158;
    assign _5 = _161;
    always @(posedge i$clock_0) begin
        if (i$clear_0)
            _85 <= _84;
        else
            if (i$enable_0)
                _85 <= _5;
    end
    assign o$total_count = _85;
    assign _162 = _79 == _76;
    assign _165 = _162 ? vdd : gnd;
    assign o$ready = _165;
    assign _171 = 1'b0;
    always @(posedge i$clock_0) begin
        if (i$clear_0)
            _170 <= _171;
        else
            if (i$enable_0)
                _170 <= o$result$last;
    end
    assign _172 = _167 ? _171 : _170;
    assign o$last_out = _172;
    assign o$last_in = _191;
    assign o$idle = _167;
    assign i$data_in$valid1 = _223;
    always @(posedge i$clock) begin
        if (i$clear)
            _226 <= _171;
        else
            if (i$enable)
                _226 <= i$data_in$valid1;
    end
    always @(posedge i$clock) begin
        if (i$clear)
            _229 <= _171;
        else
            if (i$enable)
                _229 <= _226;
    end
    always @(posedge i$clock) begin
        if (i$clear)
            _232 <= _171;
        else
            if (i$enable)
                _232 <= _229;
    end
    assign o$result$valid = _232;
    always @(posedge i$clock_0) begin
        if (i$clear_0)
            _235 <= _171;
        else
            if (i$enable_0)
                _235 <= o$result$valid;
    end
    assign _237 = _167 ? _171 : _235;
    assign o$data_out_valid = _237;
    assign _1013 = 4'b0100;
    assign _1008 = _982[0:0];
    assign _1007 = 3'b000;
    assign _1009 = { _1007,
                     _1008 };
    assign _1005 = _982[1:1];
    assign _1006 = { _1007,
                     _1005 };
    assign _1010 = _1006 + _1009;
    assign _1001 = _982[2:2];
    assign _1002 = { _1007,
                     _1001 };
    assign _998 = _982[3:3];
    assign _999 = { _1007,
                    _998 };
    assign _1003 = _999 + _1002;
    assign _1011 = _1003 + _1010;
    assign _993 = _982[4:4];
    assign _994 = { _1007,
                    _993 };
    assign _990 = _982[5:5];
    assign _991 = { _1007,
                    _990 };
    assign _995 = _991 + _994;
    assign _986 = _982[6:6];
    assign _987 = { _1007,
                    _986 };
    assign _981 = _350[0:0];
    assign _980 = _345[0:0];
    assign _979 = _343[0:0];
    assign _978 = _316[0:0];
    assign _977 = _311[0:0];
    assign _976 = _300[0:0];
    assign _975 = _295[0:0];
    assign _974 = _293[0:0];
    assign _982 = { _974,
                    _975,
                    _976,
                    _977,
                    _978,
                    _979,
                    _980,
                    _981 };
    assign _983 = _982[7:7];
    assign _984 = { _1007,
                    _983 };
    assign _988 = _984 + _987;
    assign _996 = _988 + _995;
    assign _1012 = _996 + _1011;
    assign _1014 = _1012 < _1013;
    assign _966 = _940[0:0];
    assign _967 = { _1007,
                    _966 };
    assign _963 = _940[1:1];
    assign _964 = { _1007,
                    _963 };
    assign _968 = _964 + _967;
    assign _959 = _940[2:2];
    assign _960 = { _1007,
                    _959 };
    assign _956 = _940[3:3];
    assign _957 = { _1007,
                    _956 };
    assign _961 = _957 + _960;
    assign _969 = _961 + _968;
    assign _951 = _940[4:4];
    assign _952 = { _1007,
                    _951 };
    assign _948 = _940[5:5];
    assign _949 = { _1007,
                    _948 };
    assign _953 = _949 + _952;
    assign _944 = _940[6:6];
    assign _945 = { _1007,
                    _944 };
    assign _939 = _350[1:1];
    assign _938 = _345[1:1];
    assign _937 = _343[1:1];
    assign _936 = _316[1:1];
    assign _935 = _311[1:1];
    assign _934 = _300[1:1];
    assign _933 = _295[1:1];
    assign _932 = _293[1:1];
    assign _940 = { _932,
                    _933,
                    _934,
                    _935,
                    _936,
                    _937,
                    _938,
                    _939 };
    assign _941 = _940[7:7];
    assign _942 = { _1007,
                    _941 };
    assign _946 = _942 + _945;
    assign _954 = _946 + _953;
    assign _970 = _954 + _969;
    assign _972 = _970 < _1013;
    assign _924 = _898[0:0];
    assign _925 = { _1007,
                    _924 };
    assign _921 = _898[1:1];
    assign _922 = { _1007,
                    _921 };
    assign _926 = _922 + _925;
    assign _917 = _898[2:2];
    assign _918 = { _1007,
                    _917 };
    assign _914 = _898[3:3];
    assign _915 = { _1007,
                    _914 };
    assign _919 = _915 + _918;
    assign _927 = _919 + _926;
    assign _909 = _898[4:4];
    assign _910 = { _1007,
                    _909 };
    assign _906 = _898[5:5];
    assign _907 = { _1007,
                    _906 };
    assign _911 = _907 + _910;
    assign _902 = _898[6:6];
    assign _903 = { _1007,
                    _902 };
    assign _897 = _350[2:2];
    assign _896 = _345[2:2];
    assign _895 = _343[2:2];
    assign _894 = _316[2:2];
    assign _893 = _311[2:2];
    assign _892 = _300[2:2];
    assign _891 = _295[2:2];
    assign _890 = _293[2:2];
    assign _898 = { _890,
                    _891,
                    _892,
                    _893,
                    _894,
                    _895,
                    _896,
                    _897 };
    assign _899 = _898[7:7];
    assign _900 = { _1007,
                    _899 };
    assign _904 = _900 + _903;
    assign _912 = _904 + _911;
    assign _928 = _912 + _927;
    assign _930 = _928 < _1013;
    assign _882 = _856[0:0];
    assign _883 = { _1007,
                    _882 };
    assign _879 = _856[1:1];
    assign _880 = { _1007,
                    _879 };
    assign _884 = _880 + _883;
    assign _875 = _856[2:2];
    assign _876 = { _1007,
                    _875 };
    assign _872 = _856[3:3];
    assign _873 = { _1007,
                    _872 };
    assign _877 = _873 + _876;
    assign _885 = _877 + _884;
    assign _867 = _856[4:4];
    assign _868 = { _1007,
                    _867 };
    assign _864 = _856[5:5];
    assign _865 = { _1007,
                    _864 };
    assign _869 = _865 + _868;
    assign _860 = _856[6:6];
    assign _861 = { _1007,
                    _860 };
    assign _855 = _350[3:3];
    assign _854 = _345[3:3];
    assign _853 = _343[3:3];
    assign _852 = _316[3:3];
    assign _851 = _311[3:3];
    assign _850 = _300[3:3];
    assign _849 = _295[3:3];
    assign _848 = _293[3:3];
    assign _856 = { _848,
                    _849,
                    _850,
                    _851,
                    _852,
                    _853,
                    _854,
                    _855 };
    assign _857 = _856[7:7];
    assign _858 = { _1007,
                    _857 };
    assign _862 = _858 + _861;
    assign _870 = _862 + _869;
    assign _886 = _870 + _885;
    assign _888 = _886 < _1013;
    assign _840 = _814[0:0];
    assign _841 = { _1007,
                    _840 };
    assign _837 = _814[1:1];
    assign _838 = { _1007,
                    _837 };
    assign _842 = _838 + _841;
    assign _833 = _814[2:2];
    assign _834 = { _1007,
                    _833 };
    assign _830 = _814[3:3];
    assign _831 = { _1007,
                    _830 };
    assign _835 = _831 + _834;
    assign _843 = _835 + _842;
    assign _825 = _814[4:4];
    assign _826 = { _1007,
                    _825 };
    assign _822 = _814[5:5];
    assign _823 = { _1007,
                    _822 };
    assign _827 = _823 + _826;
    assign _818 = _814[6:6];
    assign _819 = { _1007,
                    _818 };
    assign _813 = _350[4:4];
    assign _812 = _345[4:4];
    assign _811 = _343[4:4];
    assign _810 = _316[4:4];
    assign _809 = _311[4:4];
    assign _808 = _300[4:4];
    assign _807 = _295[4:4];
    assign _806 = _293[4:4];
    assign _814 = { _806,
                    _807,
                    _808,
                    _809,
                    _810,
                    _811,
                    _812,
                    _813 };
    assign _815 = _814[7:7];
    assign _816 = { _1007,
                    _815 };
    assign _820 = _816 + _819;
    assign _828 = _820 + _827;
    assign _844 = _828 + _843;
    assign _846 = _844 < _1013;
    assign _798 = _772[0:0];
    assign _799 = { _1007,
                    _798 };
    assign _795 = _772[1:1];
    assign _796 = { _1007,
                    _795 };
    assign _800 = _796 + _799;
    assign _791 = _772[2:2];
    assign _792 = { _1007,
                    _791 };
    assign _788 = _772[3:3];
    assign _789 = { _1007,
                    _788 };
    assign _793 = _789 + _792;
    assign _801 = _793 + _800;
    assign _783 = _772[4:4];
    assign _784 = { _1007,
                    _783 };
    assign _780 = _772[5:5];
    assign _781 = { _1007,
                    _780 };
    assign _785 = _781 + _784;
    assign _776 = _772[6:6];
    assign _777 = { _1007,
                    _776 };
    assign _771 = _350[5:5];
    assign _770 = _345[5:5];
    assign _769 = _343[5:5];
    assign _768 = _316[5:5];
    assign _767 = _311[5:5];
    assign _766 = _300[5:5];
    assign _765 = _295[5:5];
    assign _764 = _293[5:5];
    assign _772 = { _764,
                    _765,
                    _766,
                    _767,
                    _768,
                    _769,
                    _770,
                    _771 };
    assign _773 = _772[7:7];
    assign _774 = { _1007,
                    _773 };
    assign _778 = _774 + _777;
    assign _786 = _778 + _785;
    assign _802 = _786 + _801;
    assign _804 = _802 < _1013;
    assign _756 = _730[0:0];
    assign _757 = { _1007,
                    _756 };
    assign _753 = _730[1:1];
    assign _754 = { _1007,
                    _753 };
    assign _758 = _754 + _757;
    assign _749 = _730[2:2];
    assign _750 = { _1007,
                    _749 };
    assign _746 = _730[3:3];
    assign _747 = { _1007,
                    _746 };
    assign _751 = _747 + _750;
    assign _759 = _751 + _758;
    assign _741 = _730[4:4];
    assign _742 = { _1007,
                    _741 };
    assign _738 = _730[5:5];
    assign _739 = { _1007,
                    _738 };
    assign _743 = _739 + _742;
    assign _734 = _730[6:6];
    assign _735 = { _1007,
                    _734 };
    assign _729 = _350[6:6];
    assign _728 = _345[6:6];
    assign _727 = _343[6:6];
    assign _726 = _316[6:6];
    assign _725 = _311[6:6];
    assign _724 = _300[6:6];
    assign _723 = _295[6:6];
    assign _722 = _293[6:6];
    assign _730 = { _722,
                    _723,
                    _724,
                    _725,
                    _726,
                    _727,
                    _728,
                    _729 };
    assign _731 = _730[7:7];
    assign _732 = { _1007,
                    _731 };
    assign _736 = _732 + _735;
    assign _744 = _736 + _743;
    assign _760 = _744 + _759;
    assign _762 = _760 < _1013;
    assign _714 = _688[0:0];
    assign _715 = { _1007,
                    _714 };
    assign _711 = _688[1:1];
    assign _712 = { _1007,
                    _711 };
    assign _716 = _712 + _715;
    assign _707 = _688[2:2];
    assign _708 = { _1007,
                    _707 };
    assign _704 = _688[3:3];
    assign _705 = { _1007,
                    _704 };
    assign _709 = _705 + _708;
    assign _717 = _709 + _716;
    assign _699 = _688[4:4];
    assign _700 = { _1007,
                    _699 };
    assign _696 = _688[5:5];
    assign _697 = { _1007,
                    _696 };
    assign _701 = _697 + _700;
    assign _692 = _688[6:6];
    assign _693 = { _1007,
                    _692 };
    assign _687 = _350[7:7];
    assign _686 = _345[7:7];
    assign _685 = _343[7:7];
    assign _684 = _316[7:7];
    assign _683 = _311[7:7];
    assign _682 = _300[7:7];
    assign _681 = _295[7:7];
    assign _680 = _293[7:7];
    assign _688 = { _680,
                    _681,
                    _682,
                    _683,
                    _684,
                    _685,
                    _686,
                    _687 };
    assign _689 = _688[7:7];
    assign _690 = { _1007,
                    _689 };
    assign _694 = _690 + _693;
    assign _702 = _694 + _701;
    assign _718 = _702 + _717;
    assign _720 = _718 < _1013;
    assign _672 = _646[0:0];
    assign _673 = { _1007,
                    _672 };
    assign _669 = _646[1:1];
    assign _670 = { _1007,
                    _669 };
    assign _674 = _670 + _673;
    assign _665 = _646[2:2];
    assign _666 = { _1007,
                    _665 };
    assign _662 = _646[3:3];
    assign _663 = { _1007,
                    _662 };
    assign _667 = _663 + _666;
    assign _675 = _667 + _674;
    assign _657 = _646[4:4];
    assign _658 = { _1007,
                    _657 };
    assign _654 = _646[5:5];
    assign _655 = { _1007,
                    _654 };
    assign _659 = _655 + _658;
    assign _650 = _646[6:6];
    assign _651 = { _1007,
                    _650 };
    assign _645 = _350[8:8];
    assign _644 = _345[8:8];
    assign _643 = _343[8:8];
    assign _642 = _316[8:8];
    assign _641 = _311[8:8];
    assign _640 = _300[8:8];
    assign _639 = _295[8:8];
    assign _638 = _293[8:8];
    assign _646 = { _638,
                    _639,
                    _640,
                    _641,
                    _642,
                    _643,
                    _644,
                    _645 };
    assign _647 = _646[7:7];
    assign _648 = { _1007,
                    _647 };
    assign _652 = _648 + _651;
    assign _660 = _652 + _659;
    assign _676 = _660 + _675;
    assign _678 = _676 < _1013;
    assign _630 = _604[0:0];
    assign _631 = { _1007,
                    _630 };
    assign _627 = _604[1:1];
    assign _628 = { _1007,
                    _627 };
    assign _632 = _628 + _631;
    assign _623 = _604[2:2];
    assign _624 = { _1007,
                    _623 };
    assign _620 = _604[3:3];
    assign _621 = { _1007,
                    _620 };
    assign _625 = _621 + _624;
    assign _633 = _625 + _632;
    assign _615 = _604[4:4];
    assign _616 = { _1007,
                    _615 };
    assign _612 = _604[5:5];
    assign _613 = { _1007,
                    _612 };
    assign _617 = _613 + _616;
    assign _608 = _604[6:6];
    assign _609 = { _1007,
                    _608 };
    assign _603 = _350[9:9];
    assign _602 = _345[9:9];
    assign _601 = _343[9:9];
    assign _600 = _316[9:9];
    assign _599 = _311[9:9];
    assign _598 = _300[9:9];
    assign _597 = _295[9:9];
    assign _596 = _293[9:9];
    assign _604 = { _596,
                    _597,
                    _598,
                    _599,
                    _600,
                    _601,
                    _602,
                    _603 };
    assign _605 = _604[7:7];
    assign _606 = { _1007,
                    _605 };
    assign _610 = _606 + _609;
    assign _618 = _610 + _617;
    assign _634 = _618 + _633;
    assign _636 = _634 < _1013;
    assign _588 = _562[0:0];
    assign _589 = { _1007,
                    _588 };
    assign _585 = _562[1:1];
    assign _586 = { _1007,
                    _585 };
    assign _590 = _586 + _589;
    assign _581 = _562[2:2];
    assign _582 = { _1007,
                    _581 };
    assign _578 = _562[3:3];
    assign _579 = { _1007,
                    _578 };
    assign _583 = _579 + _582;
    assign _591 = _583 + _590;
    assign _573 = _562[4:4];
    assign _574 = { _1007,
                    _573 };
    assign _570 = _562[5:5];
    assign _571 = { _1007,
                    _570 };
    assign _575 = _571 + _574;
    assign _566 = _562[6:6];
    assign _567 = { _1007,
                    _566 };
    assign _561 = _350[10:10];
    assign _560 = _345[10:10];
    assign _559 = _343[10:10];
    assign _558 = _316[10:10];
    assign _557 = _311[10:10];
    assign _556 = _300[10:10];
    assign _555 = _295[10:10];
    assign _554 = _293[10:10];
    assign _562 = { _554,
                    _555,
                    _556,
                    _557,
                    _558,
                    _559,
                    _560,
                    _561 };
    assign _563 = _562[7:7];
    assign _564 = { _1007,
                    _563 };
    assign _568 = _564 + _567;
    assign _576 = _568 + _575;
    assign _592 = _576 + _591;
    assign _594 = _592 < _1013;
    assign _546 = _520[0:0];
    assign _547 = { _1007,
                    _546 };
    assign _543 = _520[1:1];
    assign _544 = { _1007,
                    _543 };
    assign _548 = _544 + _547;
    assign _539 = _520[2:2];
    assign _540 = { _1007,
                    _539 };
    assign _536 = _520[3:3];
    assign _537 = { _1007,
                    _536 };
    assign _541 = _537 + _540;
    assign _549 = _541 + _548;
    assign _531 = _520[4:4];
    assign _532 = { _1007,
                    _531 };
    assign _528 = _520[5:5];
    assign _529 = { _1007,
                    _528 };
    assign _533 = _529 + _532;
    assign _524 = _520[6:6];
    assign _525 = { _1007,
                    _524 };
    assign _519 = _350[11:11];
    assign _518 = _345[11:11];
    assign _517 = _343[11:11];
    assign _516 = _316[11:11];
    assign _515 = _311[11:11];
    assign _514 = _300[11:11];
    assign _513 = _295[11:11];
    assign _512 = _293[11:11];
    assign _520 = { _512,
                    _513,
                    _514,
                    _515,
                    _516,
                    _517,
                    _518,
                    _519 };
    assign _521 = _520[7:7];
    assign _522 = { _1007,
                    _521 };
    assign _526 = _522 + _525;
    assign _534 = _526 + _533;
    assign _550 = _534 + _549;
    assign _552 = _550 < _1013;
    assign _504 = _478[0:0];
    assign _505 = { _1007,
                    _504 };
    assign _501 = _478[1:1];
    assign _502 = { _1007,
                    _501 };
    assign _506 = _502 + _505;
    assign _497 = _478[2:2];
    assign _498 = { _1007,
                    _497 };
    assign _494 = _478[3:3];
    assign _495 = { _1007,
                    _494 };
    assign _499 = _495 + _498;
    assign _507 = _499 + _506;
    assign _489 = _478[4:4];
    assign _490 = { _1007,
                    _489 };
    assign _486 = _478[5:5];
    assign _487 = { _1007,
                    _486 };
    assign _491 = _487 + _490;
    assign _482 = _478[6:6];
    assign _483 = { _1007,
                    _482 };
    assign _477 = _350[12:12];
    assign _476 = _345[12:12];
    assign _475 = _343[12:12];
    assign _474 = _316[12:12];
    assign _473 = _311[12:12];
    assign _472 = _300[12:12];
    assign _471 = _295[12:12];
    assign _470 = _293[12:12];
    assign _478 = { _470,
                    _471,
                    _472,
                    _473,
                    _474,
                    _475,
                    _476,
                    _477 };
    assign _479 = _478[7:7];
    assign _480 = { _1007,
                    _479 };
    assign _484 = _480 + _483;
    assign _492 = _484 + _491;
    assign _508 = _492 + _507;
    assign _510 = _508 < _1013;
    assign _462 = _436[0:0];
    assign _463 = { _1007,
                    _462 };
    assign _459 = _436[1:1];
    assign _460 = { _1007,
                    _459 };
    assign _464 = _460 + _463;
    assign _455 = _436[2:2];
    assign _456 = { _1007,
                    _455 };
    assign _452 = _436[3:3];
    assign _453 = { _1007,
                    _452 };
    assign _457 = _453 + _456;
    assign _465 = _457 + _464;
    assign _447 = _436[4:4];
    assign _448 = { _1007,
                    _447 };
    assign _444 = _436[5:5];
    assign _445 = { _1007,
                    _444 };
    assign _449 = _445 + _448;
    assign _440 = _436[6:6];
    assign _441 = { _1007,
                    _440 };
    assign _435 = _350[13:13];
    assign _434 = _345[13:13];
    assign _433 = _343[13:13];
    assign _432 = _316[13:13];
    assign _431 = _311[13:13];
    assign _430 = _300[13:13];
    assign _429 = _295[13:13];
    assign _428 = _293[13:13];
    assign _436 = { _428,
                    _429,
                    _430,
                    _431,
                    _432,
                    _433,
                    _434,
                    _435 };
    assign _437 = _436[7:7];
    assign _438 = { _1007,
                    _437 };
    assign _442 = _438 + _441;
    assign _450 = _442 + _449;
    assign _466 = _450 + _465;
    assign _468 = _466 < _1013;
    assign _420 = _394[0:0];
    assign _421 = { _1007,
                    _420 };
    assign _417 = _394[1:1];
    assign _418 = { _1007,
                    _417 };
    assign _422 = _418 + _421;
    assign _413 = _394[2:2];
    assign _414 = { _1007,
                    _413 };
    assign _410 = _394[3:3];
    assign _411 = { _1007,
                    _410 };
    assign _415 = _411 + _414;
    assign _423 = _415 + _422;
    assign _405 = _394[4:4];
    assign _406 = { _1007,
                    _405 };
    assign _402 = _394[5:5];
    assign _403 = { _1007,
                    _402 };
    assign _407 = _403 + _406;
    assign _398 = _394[6:6];
    assign _399 = { _1007,
                    _398 };
    assign _393 = _350[14:14];
    assign _392 = _345[14:14];
    assign _391 = _343[14:14];
    assign _390 = _316[14:14];
    assign _389 = _311[14:14];
    assign _388 = _300[14:14];
    assign _387 = _295[14:14];
    assign _386 = _293[14:14];
    assign _394 = { _386,
                    _387,
                    _388,
                    _389,
                    _390,
                    _391,
                    _392,
                    _393 };
    assign _395 = _394[7:7];
    assign _396 = { _1007,
                    _395 };
    assign _400 = _396 + _399;
    assign _408 = _400 + _407;
    assign _424 = _408 + _423;
    assign _426 = _424 < _1013;
    assign _378 = _352[0:0];
    assign _379 = { _1007,
                    _378 };
    assign _375 = _352[1:1];
    assign _376 = { _1007,
                    _375 };
    assign _380 = _376 + _379;
    assign _371 = _352[2:2];
    assign _372 = { _1007,
                    _371 };
    assign _368 = _352[3:3];
    assign _369 = { _1007,
                    _368 };
    assign _373 = _369 + _372;
    assign _381 = _373 + _380;
    assign _363 = _352[4:4];
    assign _364 = { _1007,
                    _363 };
    assign _360 = _352[5:5];
    assign _361 = { _1007,
                    _360 };
    assign _365 = _361 + _364;
    assign _356 = _352[6:6];
    assign _357 = { _1007,
                    _356 };
    assign _347 = _340[46:0];
    assign _349 = { _347,
                    _171 };
    assign _350 = _349[31:16];
    assign _351 = _350[15:15];
    assign _345 = _340[31:16];
    assign _346 = _345[15:15];
    assign _338 = _325 & _287;
    assign _339 = _338 & _329;
    assign _337 = _325 & _332;
    assign i$data_in$d2 = i$data_in;
    always @(posedge i$clock) begin
        if (i$clear)
            _329 <= _72;
        else
            if (i$enable)
                _329 <= i$data_in$d2;
    end
    always @(posedge i$clock) begin
        if (i$clear)
            _332 <= _72;
        else
            if (i$enable)
                _332 <= _329;
    end
    always @(posedge i$clock) begin
        if (i$clear)
            _335 <= _72;
        else
            if (i$enable)
                _335 <= _332;
    end
    assign i$data_in$bottom1 = _238;
    always @(posedge i$clock) begin
        if (i$clear)
            _321 <= _171;
        else
            if (i$enable)
                _321 <= i$data_in$bottom1;
    end
    always @(posedge i$clock) begin
        if (i$clear)
            _324 <= _171;
        else
            if (i$enable)
                _324 <= _321;
    end
    assign _325 = _324 ? _72 : _259;
    assign _326 = _325 & _268;
    assign _336 = _326 & _335;
    assign _340 = { _336,
                    _337,
                    _339 };
    assign _341 = _340[47:1];
    assign _342 = { _171,
                    _341 };
    assign _343 = _342[31:16];
    assign _344 = _343[15:15];
    assign _313 = _308[46:0];
    assign _315 = { _313,
                    _171 };
    assign _316 = _315[31:16];
    assign _317 = _316[15:15];
    assign _307 = _287 & _67;
    always @(posedge i$clock) begin
        if (i$clear)
            _305 <= _72;
        else
            if (i$enable)
                _305 <= _70;
    end
    assign _306 = _268 & _305;
    assign _308 = { _306,
                    _70,
                    _307 };
    assign _309 = _308[47:1];
    assign _310 = { _171,
                    _309 };
    assign _311 = _310[31:16];
    assign _312 = _311[15:15];
    assign _297 = _290[46:0];
    assign _299 = { _297,
                    _171 };
    assign _300 = _299[31:16];
    assign _301 = _300[15:15];
    assign _295 = _290[31:16];
    assign _296 = _295[15:15];
    assign i$data_in$right1 = _239;
    always @(posedge i$clock) begin
        if (i$clear)
            _283 <= _171;
        else
            if (i$enable)
                _283 <= i$data_in$right1;
    end
    always @(posedge i$clock) begin
        if (i$clear)
            _286 <= _171;
        else
            if (i$enable)
                _286 <= _283;
    end
    assign _287 = _286 ? _72 : _259;
    assign _288 = _261 & _287;
    assign _289 = _288 & _272;
    assign _280 = _261 & _275;
    assign _223 = _222[17:17];
    assign _238 = _222[19:19];
    assign _239 = _222[21:21];
    assign _247 = { _239,
                    _243,
                    _238,
                    _244,
                    _223,
                    _245,
                    _246 };
    always @(posedge i$clock_0) begin
        if (_220)
            _248[_184] <= _247;
    end
    assign _241 = 10'b0000000000;
    always @(posedge i$clock_0) begin
        if (_204)
            _242 <= _198;
    end
    assign _249 = _248[_242];
    assign _250 = _249[15:0];
    assign i$data_in$d0 = _250;
    always @(posedge i$clock) begin
        if (i$clear)
            _272 <= _72;
        else
            if (i$enable)
                _272 <= i$data_in$d0;
    end
    always @(posedge i$clock) begin
        if (i$clear)
            _275 <= _72;
        else
            if (i$enable)
                _275 <= _272;
    end
    always @(posedge i$clock) begin
        if (i$clear)
            _278 <= _72;
        else
            if (i$enable)
                _278 <= _275;
    end
    assign _243 = _222[20:20];
    assign i$data_in$left1 = _243;
    always @(posedge i$clock) begin
        if (i$clear)
            _264 <= _171;
        else
            if (i$enable)
                _264 <= i$data_in$left1;
    end
    always @(posedge i$clock) begin
        if (i$clear)
            _267 <= _171;
        else
            if (i$enable)
                _267 <= _264;
    end
    assign _268 = _267 ? _72 : _259;
    assign _259 = 16'b1111111111111111;
    assign _244 = _222[18:18];
    assign i$data_in$top1 = _244;
    always @(posedge i$clock) begin
        if (i$clear)
            _255 <= _171;
        else
            if (i$enable)
                _255 <= i$data_in$top1;
    end
    always @(posedge i$clock) begin
        if (i$clear)
            _258 <= _171;
        else
            if (i$enable)
                _258 <= _255;
    end
    assign _261 = _258 ? _72 : _259;
    assign _269 = _261 & _268;
    assign _279 = _269 & _278;
    assign _290 = { _279,
                    _280,
                    _289 };
    assign _291 = _290[47:1];
    assign _292 = { _171,
                    _291 };
    assign _293 = _292[31:16];
    assign _294 = _293[15:15];
    assign _352 = { _294,
                    _296,
                    _301,
                    _312,
                    _317,
                    _344,
                    _346,
                    _351 };
    assign _353 = _352[7:7];
    assign _354 = { _1007,
                    _353 };
    assign _358 = _354 + _357;
    assign _366 = _358 + _365;
    assign _382 = _366 + _381;
    assign _384 = _382 < _1013;
    assign _1015 = { _384,
                     _426,
                     _468,
                     _510,
                     _552,
                     _594,
                     _636,
                     _678,
                     _720,
                     _762,
                     _804,
                     _846,
                     _888,
                     _930,
                     _972,
                     _1014 };
    assign _1016 = ~ _1015;
    assign _246 = _222[15:0];
    assign i$data_in$d1 = _246;
    always @(posedge i$clock) begin
        if (i$clear)
            _67 <= _72;
        else
            if (i$enable)
                _67 <= i$data_in$d1;
    end
    always @(posedge i$clock) begin
        if (i$clear)
            _70 <= _72;
        else
            if (i$enable)
                _70 <= _67;
    end
    assign _1017 = _70 & _1016;
    always @(posedge i$clock) begin
        if (i$clear)
            _1020 <= _72;
        else
            if (i$enable)
                _1020 <= _1017;
    end
    assign o$result$d = _1020;
    always @(posedge i$clock_0) begin
        if (i$clear_0)
            _1079 <= _72;
        else
            if (i$enable_0)
                _1079 <= o$result$d;
    end
    assign vdd = 1'b1;
    assign gnd = 1'b0;
    assign _75 = 2'b00;
    assign _1075 = i$start ? _79 : _76;
    assign _1072 = _191 ? _81 : _76;
    assign _1073 = i$data_in_valid ? _1072 : _76;
    assign i$enable = i$enable_0;
    assign i$clear = i$clear_0;
    assign i$clock = i$clock_0;
    assign _218 = _81 == _76;
    assign _217 = _79 == _76;
    assign _219 = _217 | _218;
    assign _220 = i$enable_0 & _219;
    assign _32 = data_in;
    assign i$data_in = _32;
    assign _185 = 10'b0000000001;
    assign _186 = _184 + _185;
    assign _190 = _186 == _189;
    assign _177 = _175 + _185;
    assign _181 = _177 == _180;
    assign _191 = _181 & _190;
    assign _215 = _175 == _241;
    assign _35 = row_size;
    assign i$row_size = _35;
    assign _1022 = i$start ? i$row_size : _180;
    assign _1021 = _76 == _75;
    assign _1023 = _1021 ? _1022 : _180;
    assign _37 = _1023;
    always @(posedge i$clock_0) begin
        if (i$clear_0)
            _180 <= _241;
        else
            if (i$enable_0)
                _180 <= _37;
    end
    assign _1038 = i$start ? _241 : _175;
    assign _1034 = _1029 ? _1031 : _175;
    assign _1035 = i$data_in_valid ? _1034 : _175;
    assign _1031 = _175 + _185;
    assign _1032 = _1029 ? _1031 : _175;
    assign _1026 = _76 == _81;
    assign _1033 = _1026 ? _1032 : _175;
    assign _1025 = _76 == _79;
    assign _1036 = _1025 ? _1035 : _1033;
    assign _1024 = _76 == _75;
    assign _1039 = _1024 ? _1038 : _1036;
    assign _38 = _1039;
    always @(posedge i$clock_0) begin
        if (i$clear_0)
            _175 <= _241;
        else
            if (i$enable_0)
                _175 <= _38;
    end
    assign _212 = _175 + _185;
    assign _213 = _212 == _180;
    assign _210 = _184 == _241;
    assign _207 = _184 + _185;
    assign _208 = _207 == _189;
    assign _216 = { _208,
                    _210,
                    _213,
                    _215,
                    i$data_in_valid,
                    _191,
                    i$data_in };
    always @(posedge i$clock_0) begin
        if (_220)
            _221[_184] <= _216;
    end
    assign _202 = _81 == _76;
    assign _201 = _79 == _76;
    assign _203 = _201 | _202;
    assign _204 = i$enable_0 & _203;
    assign _197 = _184 + _185;
    assign _1053 = i$start ? _241 : _184;
    assign _1049 = _1029 ? _241 : _1028;
    assign _40 = data_in_valid;
    assign i$data_in_valid = _40;
    assign _1050 = i$data_in_valid ? _1049 : _184;
    assign _43 = enable;
    assign i$enable_0 = _43;
    assign _46 = clear;
    assign i$clear_0 = _46;
    assign _49 = clock;
    assign i$clock_0 = _49;
    assign _52 = col_size;
    assign i$col_size = _52;
    assign _55 = start;
    assign i$start = _55;
    assign _1041 = i$start ? i$col_size : _189;
    assign _1040 = _76 == _75;
    assign _1042 = _1040 ? _1041 : _189;
    assign _57 = _1042;
    always @(posedge i$clock_0) begin
        if (i$clear_0)
            _189 <= _241;
        else
            if (i$enable_0)
                _189 <= _57;
    end
    assign _1028 = _184 + _185;
    assign _1029 = _1028 == _189;
    assign _1047 = _1029 ? _241 : _1028;
    assign _1045 = _76 == _81;
    assign _1048 = _1045 ? _1047 : _184;
    assign _1044 = _76 == _79;
    assign _1051 = _1044 ? _1050 : _1048;
    assign _1043 = _76 == _75;
    assign _1054 = _1043 ? _1053 : _1051;
    assign _58 = _1054;
    always @(posedge i$clock_0) begin
        if (i$clear_0)
            _184 <= _241;
        else
            if (i$enable_0)
                _184 <= _58;
    end
    assign _193 = _184 + _185;
    assign _194 = _193 < _189;
    assign _198 = _194 ? _197 : _241;
    always @(posedge i$clock_0) begin
        if (_204)
            _205 <= _198;
    end
    assign _222 = _221[_205];
    assign _245 = _222[16:16];
    assign i$data_in$last1 = _245;
    always @(posedge i$clock) begin
        if (i$clear)
            _1057 <= _171;
        else
            if (i$enable)
                _1057 <= i$data_in$last1;
    end
    always @(posedge i$clock) begin
        if (i$clear)
            _1060 <= _171;
        else
            if (i$enable)
                _1060 <= _1057;
    end
    always @(posedge i$clock) begin
        if (i$clear)
            _1063 <= _171;
        else
            if (i$enable)
                _1063 <= _1060;
    end
    assign o$result$last = _1063;
    assign _61 = o$result$last;
    assign _1070 = _61 ? _1067 : _76;
    assign _1067 = 2'b11;
    assign _1068 = _76 == _1067;
    assign _1069 = _1068 ? _75 : _76;
    assign _81 = 2'b10;
    assign _1066 = _76 == _81;
    assign _1071 = _1066 ? _1070 : _1069;
    assign _79 = 2'b01;
    assign _1065 = _76 == _79;
    assign _1074 = _1065 ? _1073 : _1071;
    assign _1064 = _76 == _75;
    assign _1076 = _1064 ? _1075 : _1074;
    assign _62 = _1076;
    always @(posedge i$clock_0) begin
        if (i$clear_0)
            _76 <= _75;
        else
            if (i$enable_0)
                _76 <= _62;
    end
    assign _166 = _75 == _76;
    assign _167 = _166 ? vdd : gnd;
    assign _1081 = _167 ? _72 : _1079;
    assign o$data_out = _1081;
    assign data_out = o$data_out;
    assign data_out_valid = o$data_out_valid;
    assign idle = o$idle;
    assign last_in = o$last_in;
    assign last_out = o$last_out;
    assign ready = o$ready;
    assign total_count = o$total_count;

endmodule
